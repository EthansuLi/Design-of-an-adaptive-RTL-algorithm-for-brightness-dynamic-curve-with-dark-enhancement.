module c_tab(
	input 			clk,
	input [7:0]		idata,
	
	output reg [7:0]   	o_data // 0~255
);

always@(*) begin
	case(idata)
		0	:	o_data	<=	0	;
1	:	o_data	=	2	;
2	:	o_data	=	4	;
3	:	o_data	=	7	;
4	:	o_data	=	9	;
5	:	o_data	=	12	;
6	:	o_data	=	14	;
7	:	o_data	=	16	;
8	:	o_data	=	18	;
9	:	o_data	=	21	;
10	:	o_data	=	23	;
11	:	o_data	=	25	;
12	:	o_data	=	27	;
13	:	o_data	=	29	;
14	:	o_data	=	31	;
15	:	o_data	=	33	;
16	:	o_data	=	35	;
17	:	o_data	=	37	;
18	:	o_data	=	39	;
19	:	o_data	=	41	;
20	:	o_data	=	43	;
21	:	o_data	=	45	;
22	:	o_data	=	47	;
23	:	o_data	=	49	;
24	:	o_data	=	50	;
25	:	o_data	=	52	;
26	:	o_data	=	54	;
27	:	o_data	=	56	;
28	:	o_data	=	57	;
29	:	o_data	=	59	;
30	:	o_data	=	61	;
31	:	o_data	=	63	;
32	:	o_data	=	64	;
33	:	o_data	=	66	;
34	:	o_data	=	67	;
35	:	o_data	=	69	;
36	:	o_data	=	71	;
37	:	o_data	=	72	;
38	:	o_data	=	74	;
39	:	o_data	=	75	;
40	:	o_data	=	77	;
41	:	o_data	=	78	;
42	:	o_data	=	80	;
43	:	o_data	=	81	;
44	:	o_data	=	83	;
45	:	o_data	=	84	;
46	:	o_data	=	86	;
47	:	o_data	=	87	;
48	:	o_data	=	89	;
49	:	o_data	=	90	;
50	:	o_data	=	92	;
51	:	o_data	=	93	;
52	:	o_data	=	94	;
53	:	o_data	=	96	;
54	:	o_data	=	97	;
55	:	o_data	=	98	;
56	:	o_data	=	100	;
57	:	o_data	=	101	;
58	:	o_data	=	102	;
59	:	o_data	=	104	;
60	:	o_data	=	105	;
61	:	o_data	=	106	;
62	:	o_data	=	108	;
63	:	o_data	=	109	;
64	:	o_data	=	110	;
65	:	o_data	=	111	;
66	:	o_data	=	113	;
67	:	o_data	=	114	;
68	:	o_data	=	115	;
69	:	o_data	=	116	;
70	:	o_data	=	117	;
71	:	o_data	=	119	;
72	:	o_data	=	120	;
73	:	o_data	=	121	;
74	:	o_data	=	122	;
75	:	o_data	=	123	;
76	:	o_data	=	124	;
77	:	o_data	=	125	;
78	:	o_data	=	127	;
79	:	o_data	=	128	;
80	:	o_data	=	129	;
81	:	o_data	=	130	;
82	:	o_data	=	131	;
83	:	o_data	=	132	;
84	:	o_data	=	133	;
85	:	o_data	=	134	;
86	:	o_data	=	135	;
87	:	o_data	=	136	;
88	:	o_data	=	137	;
89	:	o_data	=	138	;
90	:	o_data	=	140	;
91	:	o_data	=	141	;
92	:	o_data	=	142	;
93	:	o_data	=	143	;
94	:	o_data	=	144	;
95	:	o_data	=	145	;
96	:	o_data	=	146	;
97	:	o_data	=	147	;
98	:	o_data	=	148	;
99	:	o_data	=	149	;
100	:	o_data	=	150	;
101	:	o_data	=	151	;
102	:	o_data	=	151	;
103	:	o_data	=	152	;
104	:	o_data	=	153	;
105	:	o_data	=	154	;
106	:	o_data	=	155	;
107	:	o_data	=	156	;
108	:	o_data	=	157	;
109	:	o_data	=	158	;
110	:	o_data	=	159	;
111	:	o_data	=	160	;
112	:	o_data	=	161	;
113	:	o_data	=	162	;
114	:	o_data	=	163	;
115	:	o_data	=	163	;
116	:	o_data	=	164	;
117	:	o_data	=	165	;
118	:	o_data	=	166	;
119	:	o_data	=	167	;
120	:	o_data	=	168	;
121	:	o_data	=	169	;
122	:	o_data	=	170	;
123	:	o_data	=	170	;
124	:	o_data	=	171	;
125	:	o_data	=	172	;
126	:	o_data	=	173	;
127	:	o_data	=	174	;
128	:	o_data	=	175	;
129	:	o_data	=	175	;
130	:	o_data	=	176	;
131	:	o_data	=	177	;
132	:	o_data	=	178	;
133	:	o_data	=	179	;
134	:	o_data	=	180	;
135	:	o_data	=	180	;
136	:	o_data	=	181	;
137	:	o_data	=	182	;
138	:	o_data	=	183	;
139	:	o_data	=	184	;
140	:	o_data	=	184	;
141	:	o_data	=	185	;
142	:	o_data	=	186	;
143	:	o_data	=	187	;
144	:	o_data	=	187	;
145	:	o_data	=	188	;
146	:	o_data	=	189	;
147	:	o_data	=	190	;
148	:	o_data	=	190	;
149	:	o_data	=	191	;
150	:	o_data	=	192	;
151	:	o_data	=	193	;
152	:	o_data	=	193	;
153	:	o_data	=	194	;
154	:	o_data	=	195	;
155	:	o_data	=	196	;
156	:	o_data	=	196	;
157	:	o_data	=	197	;
158	:	o_data	=	198	;
159	:	o_data	=	198	;
160	:	o_data	=	199	;
161	:	o_data	=	200	;
162	:	o_data	=	201	;
163	:	o_data	=	201	;
164	:	o_data	=	202	;
165	:	o_data	=	203	;
166	:	o_data	=	203	;
167	:	o_data	=	204	;
168	:	o_data	=	205	;
169	:	o_data	=	205	;
170	:	o_data	=	206	;
171	:	o_data	=	207	;
172	:	o_data	=	208	;
173	:	o_data	=	208	;
174	:	o_data	=	209	;
175	:	o_data	=	210	;
176	:	o_data	=	210	;
177	:	o_data	=	211	;
178	:	o_data	=	212	;
179	:	o_data	=	212	;
180	:	o_data	=	213	;
181	:	o_data	=	213	;
182	:	o_data	=	214	;
183	:	o_data	=	215	;
184	:	o_data	=	215	;
185	:	o_data	=	216	;
186	:	o_data	=	217	;
187	:	o_data	=	217	;
188	:	o_data	=	218	;
189	:	o_data	=	219	;
190	:	o_data	=	219	;
191	:	o_data	=	220	;
192	:	o_data	=	220	;
193	:	o_data	=	221	;
194	:	o_data	=	222	;
195	:	o_data	=	222	;
196	:	o_data	=	223	;
197	:	o_data	=	224	;
198	:	o_data	=	224	;
199	:	o_data	=	225	;
200	:	o_data	=	225	;
201	:	o_data	=	226	;
202	:	o_data	=	227	;
203	:	o_data	=	227	;
204	:	o_data	=	228	;
205	:	o_data	=	228	;
206	:	o_data	=	229	;
207	:	o_data	=	230	;
208	:	o_data	=	230	;
209	:	o_data	=	231	;
210	:	o_data	=	231	;
211	:	o_data	=	232	;
212	:	o_data	=	232	;
213	:	o_data	=	233	;
214	:	o_data	=	234	;
215	:	o_data	=	234	;
216	:	o_data	=	235	;
217	:	o_data	=	235	;
218	:	o_data	=	236	;
219	:	o_data	=	236	;
220	:	o_data	=	237	;
221	:	o_data	=	238	;
222	:	o_data	=	238	;
223	:	o_data	=	239	;
224	:	o_data	=	239	;
225	:	o_data	=	240	;
226	:	o_data	=	240	;
227	:	o_data	=	241	;
228	:	o_data	=	241	;
229	:	o_data	=	242	;
230	:	o_data	=	243	;
231	:	o_data	=	243	;
232	:	o_data	=	244	;
233	:	o_data	=	244	;
234	:	o_data	=	245	;
235	:	o_data	=	245	;
236	:	o_data	=	246	;
237	:	o_data	=	246	;
238	:	o_data	=	247	;
239	:	o_data	=	247	;
240	:	o_data	=	248	;
241	:	o_data	=	248	;
242	:	o_data	=	249	;
243	:	o_data	=	249	;
244	:	o_data	=	250	;
245	:	o_data	=	250	;
246	:	o_data	=	251	;
247	:	o_data	=	251	;
248	:	o_data	=	252	;
249	:	o_data	=	252	;
250	:	o_data	=	253	;
251	:	o_data	=	253	;
252	:	o_data	=	254	;
253	:	o_data	=	254	;
254	:	o_data	=	255	;
255	:	o_data	=	255	;
		
	default : o_data=idata;
	endcase
end

endmodule